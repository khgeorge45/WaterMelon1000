module tb;
int c = a+b;
endmodule
