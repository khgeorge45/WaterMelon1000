class monitor
endclass
